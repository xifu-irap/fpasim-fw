-- -------------------------------------------------------------------------------------------------------------
--                              Copyright (C) 2022-2030 Ken-ji de la Rosa, IRAP Toulouse.
-- -------------------------------------------------------------------------------------------------------------
--                              This file is part of the ATHENA X-IFU DRE Focal Plane Assembly simulator.
--
--                              fpasim-fw is free software: you can redistribute it and/or modify
--                              it under the terms of the GNU General Public License as published by
--                              the Free Software Foundation, either version 3 of the License, or
--                              (at your option) any later version.
--
--                              This program is distributed in the hope that it will be useful,
--                              but WITHOUT ANY WARRANTY; without even the implied warranty of
--                              MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--                              GNU General Public License for more details.
--
--                              You should have received a copy of the GNU General Public License
--                              along with this program.  If not, see <https://www.gnu.org/licenses/>.
-- -------------------------------------------------------------------------------------------------------------
--    email                   kenji.delarosa@alten.com
--    @file                   io_sync.vhd 
-- -------------------------------------------------------------------------------------------------------------
--    Automatic Generation    No
--    Code Rules Reference    SOC of design and VHDL handbook for VLSI development, CNES Edition (v2.1)
-- -------------------------------------------------------------------------------------------------------------
--    @details                
--
--    This module generates fpga specific IO component with an optional user-defined latency

--    Example0:
--      Input ports -> optionnal latency -> fpga specific IO generation -> output port
--
-- -------------------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

use work.pkg_fpasim.all;

entity io_sync is
  generic(
    g_OUTPUT_LATENCY : natural := 0  -- add latency before the output IO. Possible values: [0; max integer values[
    );
  port(

    ---------------------------------------------------------------------
    -- input
    ---------------------------------------------------------------------
    i_clk         : in  std_logic;      -- clock
    i_rst         : in  std_logic;      -- reset
    i_rst_status  : in  std_logic;      -- reset error flag(s)
    i_debug_pulse : in  std_logic;      -- error mode (transparent vs capture). Possible values: '1': delay the error(s), '0': capture the error(s)
    i_sync_valid  : in  std_logic;      -- sync valid
    i_sync        : in  std_logic;      -- sync value
    
    ---------------------------------------------------------------------
    -- output @i_out_clk
    ---------------------------------------------------------------------
    i_out_clk     : in  std_logic;  -- output clock
    -- from reset_top: @i_out_clk
    i_io_clk_rst  : in  std_logic;  -- Clock reset: Reset connected to clocking elements in the circuit
    i_io_rst      : in  std_logic;  -- Reset connected to all other elements in the circuit
    -- data
    o_sync_clk    : out std_logic;
    o_sync        : out std_logic;

    ---------------------------------------------------------------------
    -- errors/status @i_clk
    --------------------------------------------------------------------- 
    o_errors : out std_logic_vector(15 downto 0);  -- output errors
    o_status : out std_logic_vector(7 downto 0)    -- output status
    );
end entity io_sync;

architecture RTL of io_sync is


  constant c_FIFO_READ_LATENCY : natural := pkg_IO_SYNC_FIFO_READ_LATENCY;
  ---------------------------------------------------------------------
  -- FIFO
  ---------------------------------------------------------------------
  constant c_IDX0_L            : integer := 0;
  constant c_IDX0_H            : integer := c_IDX0_L + 1 - 1;

  constant c_FIFO_DEPTH : integer := 16;            --see IP
  constant c_FIFO_WIDTH : integer := c_IDX0_H + 1;  --see IP

  signal wr_rst_tmp0 : std_logic;
  signal wr_tmp0     : std_logic;
  signal data_tmp0   : std_logic_vector(c_FIFO_WIDTH - 1 downto 0);
  --signal full0        : std_logic;
  --signal wr_rst_busy0 : std_logic;

  signal errors_sync0 : std_logic_vector(3 downto 0);
  signal empty_sync0  : std_logic;

  signal rd1       : std_logic;
  signal data_tmp1 : std_logic_vector(c_FIFO_WIDTH - 1 downto 0);
  signal empty1    : std_logic;
  --signal rd_rst_busy1 : std_logic;

  signal sync_valid1 : std_logic;
  signal sync1       : std_logic;

  ---------------------------------------------------------------------
  -- optionnally add latency
  ---------------------------------------------------------------------
  signal sync_rx : std_logic;

  ---------------------------------------------------------------------
  -- oddr
  ---------------------------------------------------------------------
  signal sync_tmp : std_logic;
  signal clk_tmp  : std_logic;

  ---------------------------------------------------------------------
  -- error latching
  ---------------------------------------------------------------------
  constant NB_ERRORS_c : integer := 3;
  signal error_tmp     : std_logic_vector(NB_ERRORS_c - 1 downto 0);
  signal error_tmp_bis : std_logic_vector(NB_ERRORS_c - 1 downto 0);

begin
---------------------------------------------------------------------
  -- clock domain crossing
  ---------------------------------------------------------------------
  wr_rst_tmp0         <= i_rst;
  wr_tmp0             <= i_sync_valid;
  data_tmp0(c_IDX0_H) <= i_sync;

  inst_fifo_async_with_error : entity work.fifo_async_with_error
    generic map(
      g_CDC_SYNC_STAGES   => 2,
      g_FIFO_MEMORY_TYPE  => "auto",
      g_FIFO_READ_LATENCY => c_FIFO_READ_LATENCY,
      g_FIFO_WRITE_DEPTH  => c_FIFO_DEPTH,
      g_READ_DATA_WIDTH   => data_tmp1'length,
      g_READ_MODE         => "std",
      g_RELATED_CLOCKS    => 0,
      g_WRITE_DATA_WIDTH  => data_tmp0'length,
      ---------------------------------------------------------------------
      -- resynchronization: fifo errors/empty flag
      ---------------------------------------------------------------------
      g_SYNC_SIDE         => "wr"  -- define the clock side where status/errors is resynchronised. Possible value "wr" or "rd"

      )
    port map(
      ---------------------------------------------------------------------
      -- write side
      ---------------------------------------------------------------------
      i_wr_clk        => i_clk,
      i_wr_rst        => wr_rst_tmp0,
      i_wr_en         => wr_tmp0,
      i_wr_din        => data_tmp0,
      o_wr_full       => open,
      o_wr_rst_busy   => open,
      ---------------------------------------------------------------------
      -- read side
      ---------------------------------------------------------------------
      i_rd_clk        => i_out_clk,
      i_rd_en         => rd1,
      o_rd_dout_valid => sync_valid1,
      o_rd_dout       => data_tmp1,
      o_rd_empty      => empty1,
      o_rd_rst_busy   => open,
      ---------------------------------------------------------------------
      -- resynchronized errors/status 
      ---------------------------------------------------------------------
      o_errors_sync   => errors_sync0,
      o_empty_sync    => empty_sync0
      );

  rd1 <= '1' when empty1 = '0' else '0';

  sync1 <= data_tmp1(c_IDX0_H) and sync_valid1;


  ---------------------------------------------------------------------
  -- output: optionnally add latency before output IOs
  ---------------------------------------------------------------------
  inst_pipeliner_add_output_latency : entity work.pipeliner
    generic map(
      g_NB_PIPES   => g_OUTPUT_LATENCY,  -- number of consecutives registers. Possibles values: [0, integer max value[
      g_DATA_WIDTH => 1  -- width of the input/output data.  Possibles values: [1, integer max value[
      )
    port map(
      i_clk     => i_out_clk,           -- clock signal
      i_data(0) => sync1,               -- input data
      o_data(0) => sync_rx              -- output data with/without delay
      );

  ---------------------------------------------------------------------
  -- I/O interface
  ---------------------------------------------------------------------
  gen_io_sync : if true generate
    signal data_tmp0 : std_logic_vector(0 downto 0);
    signal data_tmp1 : std_logic_vector(0 downto 0);
  begin
    data_tmp0(0) <= sync_rx;
    inst_selectio_wiz_sync : entity work.selectio_wiz_sync
      port map(
        data_out_from_device => data_tmp0,
        data_out_to_pins     => data_tmp1,
        clk_to_pins          => clk_tmp,
        clk_in               => i_out_clk,
        clk_reset            => i_io_clk_rst,
        io_reset             => i_io_rst
        );
    sync_tmp <= data_tmp1(0);
  end generate gen_io_sync;

  ---------------------------------------------------------------------
  -- output
  ---------------------------------------------------------------------
  o_sync_clk <= clk_tmp;
  o_sync     <= sync_tmp;


  ---------------------------------------------------------------------
  -- Error latching
  ---------------------------------------------------------------------
  error_tmp(2) <= errors_sync0(2) or errors_sync0(3);  -- fifo rst error
  error_tmp(1) <= errors_sync0(1);                     -- fifo rd empty error
  error_tmp(0) <= errors_sync0(0);                     -- fifo wr full error
  gen_errors_latch : for i in error_tmp'range generate
    inst_one_error_latch : entity work.one_error_latch
      port map(
        i_clk         => i_clk,
        i_rst         => i_rst_status,
        i_debug_pulse => i_debug_pulse,
        i_error       => error_tmp(i),
        o_error       => error_tmp_bis(i)
        );
  end generate gen_errors_latch;

  o_errors(15 downto 3) <= (others => '0');
  o_errors(2)           <= error_tmp_bis(2);  -- fifo rst error
  o_errors(1)           <= error_tmp_bis(1);  -- fifo rd empty error
  o_errors(0)           <= error_tmp_bis(0);  -- fifo wr full error

  o_status(7 downto 1) <= (others => '0');
  o_status(0)          <= empty_sync0;

  ---------------------------------------------------------------------
  -- for simulation only
  ---------------------------------------------------------------------
  assert not (error_tmp_bis(2) = '1') report "[io_sync] => FIFO is used before the end of the initialization " severity error;
  assert not (error_tmp_bis(1) = '1') report "[io_sync] => FIFO read an empty FIFO" severity error;
  assert not (error_tmp_bis(0) = '1') report "[io_sync] => FIFO write a full FIFO" severity error;

end architecture RTL;
