-- -------------------------------------------------------------------------------------------------------------
--                              Copyright (C) 2022-2030 Ken-ji de la Rosa, IRAP Toulouse.
-- -------------------------------------------------------------------------------------------------------------
--                              This file is part of the ATHENA X-IFU DRE Focal Plane Assembly simulator.
--
--                              fpasim-fw is free software: you can redistribute it and/or modify
--                              it under the terms of the GNU General Public License as published by
--                              the Free Software Foundation, either version 3 of the License, or
--                              (at your option) any later version.
--
--                              This program is distributed in the hope that it will be useful,
--                              but WITHOUT ANY WARRANTY; without even the implied warranty of
--                              MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--                              GNU General Public License for more details.
--
--                              You should have received a copy of the GNU General Public License
--                              along with this program.  If not, see <https://www.gnu.org/licenses/>.
-- -------------------------------------------------------------------------------------------------------------
--    email                   kenji.delarosa@alten.com
--!   @file                   pkg_front_panel.vhd 
-- -------------------------------------------------------------------------------------------------------------
--    Automatic Generation    No
--    Code Rules Reference    SOC of design and VHDL handbook for VLSI development, CNES Edition (v2.1)
-- -------------------------------------------------------------------------------------------------------------
--!   @details                
--
--
-- -------------------------------------------------------------------------------------------------------------

library ieee;
library std;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
use IEEE.std_logic_textio.all;

use std.textio.all;

library opal_kelly_lib;
use opal_kelly_lib.parameters.all;

package pkg_front_panel is

    type t_void is (VOID);

    ------------------------------------------------------
    -- this procedure allows to wait a number of rising edge
    -- then a margin is applied, if any
    ------------------------------------------------------
    procedure wait_nb_rising_edge_plus_margin(
        signal   i_clk            : in std_logic;
        constant i_nb_rising_edge : in natural;
        constant i_margin         : in time
    );

    type t_internal_if is record
        hi_drive   : std_logic;
        hi_cmd     : std_logic_vector(2 downto 0);
        hi_busy    : std_logic;
        hi_datain  : std_logic_vector(31 downto 0);
        hi_dataout : std_logic_vector(31 downto 0);

    end record t_internal_if;


    constant DNOP                  : std_logic_vector(2 downto 0) := "000";
    constant DReset                : std_logic_vector(2 downto 0) := "001";
    constant DWires                : std_logic_vector(2 downto 0) := "010";
    constant DUpdateWireIns        : std_logic_vector(2 downto 0) := "001";
    constant DUpdateWireOuts       : std_logic_vector(2 downto 0) := "010";
    constant DTriggers             : std_logic_vector(2 downto 0) := "011";
    constant DActivateTriggerIn    : std_logic_vector(2 downto 0) := "001";
    constant DUpdateTriggerOuts    : std_logic_vector(2 downto 0) := "010";
    constant DPipes                : std_logic_vector(2 downto 0) := "100";
    constant DWriteToPipeIn        : std_logic_vector(2 downto 0) := "001";
    constant DReadFromPipeOut      : std_logic_vector(2 downto 0) := "010";
    constant DWriteToBlockPipeIn   : std_logic_vector(2 downto 0) := "011";
    constant DReadFromBlockPipeOut : std_logic_vector(2 downto 0) := "100";
    constant DRegisters            : std_logic_vector(2 downto 0) := "101";
    constant DWriteRegister        : std_logic_vector(2 downto 0) := "001";
    constant DReadRegister         : std_logic_vector(2 downto 0) := "010";
    constant DWriteRegisterSet     : std_logic_vector(2 downto 0) := "011";
    constant DReadRegisterSet      : std_logic_vector(2 downto 0) := "100";

    type PIPEIN_ARRAY is array (integer range <>) of std_logic_vector(7 downto 0);
    type PIPEOUT_ARRAY is array (integer range <>) of std_logic_vector(7 downto 0);
    type STD_ARRAY is array (integer range <>) of std_logic_vector(31 downto 0);
    type REGISTER_ARRAY is array (integer range <>) of std_logic_vector(31 downto 0);
    
    type t_front_panel_conf is record
        pipeIn           : PIPEIN_ARRAY;

        pipeOut          : PIPEOUT_ARRAY;

        WireIns          : STD_ARRAY;   -- 32x32 array storing WireIn values
        WireOuts         : STD_ARRAY;   -- 32x32 array storing WireOut values 
        Triggered        : STD_ARRAY;   -- 32x32 array storing IsTriggered values

        u32Address       : REGISTER_ARRAY;
        u32Data          : REGISTER_ARRAY;
        u32Count         : std_logic_vector(31 downto 0);
        ReadRegisterData : std_logic_vector(31 downto 0);

        PostReadyDelay   : integer;
        ReadyCheckDelay  : integer;
        BlockDelayStates : integer;

    end record t_front_panel_conf;




    -----------------------------------------------------------------------
    -- init_front_panel_conf
    -----------------------------------------------------------------------
    impure function init_front_panel_conf(
         BlockDelayStates : in integer := 5; -- REQUIRED: # of clocks between blocks of pipe data
         ReadyCheckDelay  : in integer := 5; -- REQUIRED: # of clocks before block transfer before host interface checks for ready (0-255)
         PostReadyDelay   : in integer := 5; -- REQUIRED: # of clocks after ready is asserted and check that the block transfer begins (0-255)
         pipeInSize       : in integer := 1024; -- REQUIRED: byte (must be even) length of default PipeIn; Integer 0-2^32
         pipeOutSize      : in integer := 1024; -- REQUIRED: byte (must be even) length of default PipeOut; Integer 0-2^32
         registerSetSize  : in integer := 32 -- Size of array for register set commands.
    ) return t_front_panel_conf;

    impure function init_internal_if( dummy : in integer) return t_internal_if;

    procedure okHost_driver(
        signal i_clk : in std_logic;
        signal okUH      : out STD_LOGIC_VECTOR (4  downto 0);
        signal okHU      : in STD_LOGIC_VECTOR (2  downto 0);
        signal okUHU     : inout STD_LOGIC_VECTOR (31 downto 0);
        signal internal_if : inout t_internal_if
    );

    -----------------------------------------------------------------------
    -- Available User Task and Function Calls:
    --    FrontPanelReset;              -- Always start routine with FrontPanelReset;
    --    SetWireInValue(ep, val, mask);
    --    UpdateWireIns;
    --    UpdateWireOuts;
    --    GetWireOutValue(ep);          -- returns a 16 bit SLV
    --    ActivateTriggerIn(ep, bit);   -- bit is an integer 0-15
    --    UpdateTriggerOuts;
    --    IsTriggered(ep, mask);        -- returns a BOOLEAN
    --    WriteToPipeIn(ep, length);    -- pass pipeIn array data; length is integer
    --    ReadFromPipeOut(ep, length);  -- pass data to pipeOut array; length is integer
    --    WriteToBlockPipeIn(ep, blockSize, length);   -- pass pipeIn array data; blockSize and length are integers
    --    ReadFromBlockPipeOut(ep, blockSize, length); -- pass data to pipeOut array; blockSize and length are integers
    --    WriteRegister(addr, data);  
    --    ReadRegister(addr, data);
    --    WriteRegisterSet();  
    --    ReadRegisterSet();
    --
    -- *  Pipes operate by passing arrays of data back and forth to the user's
    --    design.  If you need multiple arrays, you can create a new procedure
    --    above and connect it to a differnet array.  More information is
    --    available in Opal Kelly documentation and online support tutorial.
    ----------------------------------------------------------------------- 
    -----------------------------------------------------------------------
    -- FrontPanelReset
    -----------------------------------------------------------------------
    procedure FrontPanelReset(signal i_clk : in std_logic; variable front_panel_conf : inout t_front_panel_conf; signal internal_if : inout t_internal_if);

    -----------------------------------------------------------------------
    -- SetWireInValue
    -----------------------------------------------------------------------
    procedure SetWireInValue(
        ep                   : in std_logic_vector(7 downto 0);
        val                  : in std_logic_vector(31 downto 0);
        mask                 : in std_logic_vector(31 downto 0);
        variable front_panel_conf : inout t_front_panel_conf
    );

    -----------------------------------------------------------------------
    -- GetWireOutValue
    -----------------------------------------------------------------------
    impure function GetWireOutValue(
        ep          : std_logic_vector;
        front_panel_conf : in t_front_panel_conf) return std_logic_vector;

    -----------------------------------------------------------------------
    -- IsTriggered
    -----------------------------------------------------------------------
    impure function IsTriggered(
        ep          : std_logic_vector;
        mask        : std_logic_vector(31 downto 0);
        front_panel_conf : t_front_panel_conf
    ) return boolean;

    -----------------------------------------------------------------------
    -- UpdateWireIns
    -----------------------------------------------------------------------
    procedure UpdateWireIns(signal   i_clk   : in std_logic;
                            variable front_panel_conf : inout t_front_panel_conf;
                            signal   internal_if   : inout t_internal_if
                           );

    -----------------------------------------------------------------------
    -- UpdateWireOuts
    -----------------------------------------------------------------------
    procedure UpdateWireOuts(
        signal   i_clk   : in std_logic;
        variable front_panel_conf : inout t_front_panel_conf;
        signal   internal_if   : inout t_internal_if
    );

    -----------------------------------------------------------------------
    -- ActivateTriggerIn
    -----------------------------------------------------------------------
    procedure ActivateTriggerIn(
        signal i_clk : in std_logic;
        ep               : in std_logic_vector(7 downto 0);
        bit              : in integer;
        signal internal_if : inout t_internal_if);

    -----------------------------------------------------------------------
    -- UpdateTriggerOuts
    -----------------------------------------------------------------------
    procedure UpdateTriggerOuts(
        signal   i_clk   : in std_logic;
        variable front_panel_conf : inout t_front_panel_conf;
        signal   internal_if   : inout t_internal_if
    );

    -----------------------------------------------------------------------
    -- WriteToPipeIn
    -----------------------------------------------------------------------
    procedure WriteToPipeIn(
        signal   i_clk   : in std_logic;
        ep                   : in std_logic_vector(7 downto 0);
        length               : in integer;
        variable front_panel_conf : inout t_front_panel_conf;
        signal   internal_if   : inout t_internal_if
    );

    -----------------------------------------------------------------------
    -- ReadFromPipeOut
    -----------------------------------------------------------------------
    procedure ReadFromPipeOut(
        signal   i_clk   : in std_logic;
        ep                   : in std_logic_vector(7 downto 0);
        length               : in integer;
        variable front_panel_conf : inout t_front_panel_conf;
        signal   internal_if   : inout t_internal_if
    );

    -----------------------------------------------------------------------
    -- WriteToBlockPipeIn
    -----------------------------------------------------------------------
    procedure WriteToBlockPipeIn(
        signal   i_clk   : in std_logic;
        ep                   : in std_logic_vector(7 downto 0);
        blockLength          : in integer;
        length               : in integer;
        variable front_panel_conf : inout t_front_panel_conf;
        signal   internal_if   : inout t_internal_if);

    -----------------------------------------------------------------------
    -- ReadFromBlockPipeOut
    -----------------------------------------------------------------------
    procedure ReadFromBlockPipeOut(
        signal   i_clk   : in std_logic;
        ep                   : in std_logic_vector(7 downto 0);
        blockLength          : in integer;
        length               : in integer;
        variable front_panel_conf : inout t_front_panel_conf;
        signal   internal_if   : inout t_internal_if);

    -----------------------------------------------------------------------
    -- WriteRegister
    -----------------------------------------------------------------------
    procedure WriteRegister(
        signal i_clk : in std_logic;
        address          : in std_logic_vector(31 downto 0);
        data             : in std_logic_vector(31 downto 0);
        signal internal_if : inout t_internal_if);

    -----------------------------------------------------------------------
    -- ReadRegister
    -----------------------------------------------------------------------
    procedure ReadRegister(
        signal i_clk : in std_logic;
        address          : in std_logic_vector(31 downto 0);
        data             : out std_logic_vector(31 downto 0);
        signal internal_if : inout t_internal_if
    );

    -----------------------------------------------------------------------
    -- WriteRegisterSet
    -----------------------------------------------------------------------
    procedure WriteRegisterSet(
        signal   i_clk   : in std_logic;
        variable front_panel_conf : inout t_front_panel_conf;
        signal   internal_if   : inout t_internal_if
    );

    -----------------------------------------------------------------------
    -- ReadRegisterSet
    -----------------------------------------------------------------------
    procedure ReadRegisterSet(
        signal   i_clk   : in std_logic;
        variable front_panel_conf : inout t_front_panel_conf;
        signal   internal_if   : inout t_internal_if);

end;

package body pkg_front_panel is

    ------------------------------------------------------
    -- this procedure allows to wait a number of rising edge
    -- then a margin is applied, if any
    ------------------------------------------------------
    procedure wait_nb_rising_edge_plus_margin(
        signal   i_clk            : in std_logic;
        constant i_nb_rising_edge : in natural;
        constant i_margin         : in time
    ) is
    begin
        -- Wait for number of rising edges
        --   if the number of rising edges = 0 => only the margin is applied, if any
        if i_nb_rising_edge /= 0 then
            for i in 1 to i_nb_rising_edge loop
                wait until rising_edge(i_clk);
            end loop;
        end if;
        -- Wait for i_margin time, if any
        wait for i_margin;
    end procedure;

    --type t_front_panel is protected body

    --variable  hi_drive   : std_logic := '0';
    --variable  hi_cmd     : std_logic_vector(2 downto 0) := "000";
    --variable  hi_busy    : std_logic;
    --variable  hi_datain  : std_logic_vector(31 downto 0) := x"00000000";
    --variable  hi_dataout : std_logic_vector(31 downto 0) := x"00000000";

    -----------------------------------------------------------------------
    -- Required data for procedures and functions
    -----------------------------------------------------------------------
    -- If you require multiple pipe arrays, you may create more arrays here
    -- duplicate the desired pipe procedures as required, change the names
    -- of the duplicated procedure to a unique identifiers, and alter the
    -- pipe array in that procedure to your newly generated arrays here.
    --type PIPEIN_ARRAY is array (0 to pipeInSize - 1) of std_logic_vector(7 downto 0);
    --variable pipeIn   : PIPEIN_ARRAY;

    --type PIPEOUT_ARRAY is array (0 to pipeOutSize - 1) of std_logic_vector(7 downto 0);
    --variable pipeOut  : PIPEOUT_ARRAY;

    --type STD_ARRAY is array (0 to 31) of std_logic_vector(31 downto 0);
    --variable WireIns    :  STD_ARRAY; -- 32x32 array storing WireIn values
    --variable WireOuts   :  STD_ARRAY; -- 32x32 array storing WireOut values 
    --variable Triggered  :  STD_ARRAY; -- 32x32 array storing IsTriggered values

    --type REGISTER_ARRAY is array (0 to registerSetSize - 1) of std_logic_vector(31 downto 0);
    --variable u32Address  : REGISTER_ARRAY;
    --variable u32Data     : REGISTER_ARRAY;
    --variable u32Count    : std_logic_vector(31 downto 0);
    --variable ReadRegisterData    : std_logic_vector(31 downto 0);

    --constant DNOP                  : std_logic_vector(2 downto 0) := "000";
    --constant DReset                : std_logic_vector(2 downto 0) := "001";
    --constant DWires                : std_logic_vector(2 downto 0) := "010";
    --constant DUpdateWireIns        : std_logic_vector(2 downto 0) := "001";
    --constant DUpdateWireOuts       : std_logic_vector(2 downto 0) := "010";
    --constant DTriggers             : std_logic_vector(2 downto 0) := "011";
    --constant DActivateTriggerIn    : std_logic_vector(2 downto 0) := "001";
    --constant DUpdateTriggerOuts    : std_logic_vector(2 downto 0) := "010";
    --constant DPipes                : std_logic_vector(2 downto 0) := "100";
    --constant DWriteToPipeIn        : std_logic_vector(2 downto 0) := "001";
    --constant DReadFromPipeOut      : std_logic_vector(2 downto 0) := "010";
    --constant DWriteToBlockPipeIn   : std_logic_vector(2 downto 0) := "011";
    --constant DReadFromBlockPipeOut : std_logic_vector(2 downto 0) := "100";
    --constant DRegisters            : std_logic_vector(2 downto 0) := "101";
    --constant DWriteRegister        : std_logic_vector(2 downto 0) := "001";
    --constant DReadRegister         : std_logic_vector(2 downto 0) := "010";
    --constant DWriteRegisterSet     : std_logic_vector(2 downto 0) := "011";
    --constant DReadRegisterSet      : std_logic_vector(2 downto 0) := "100";

    procedure okHost_driver(
        signal i_clk : in std_logic;
        signal okUH      : out STD_LOGIC_VECTOR (4  downto 0);
        signal okHU      : in STD_LOGIC_VECTOR (2  downto 0);
        signal okUHU     : inout STD_LOGIC_VECTOR (31 downto 0);
        signal internal_if : inout t_internal_if
    ) is

        --variable v_test : boolean := true;

    begin
        --while v_test = True loop
        -- okHostCalls Simulation okHostCall<->okHost Mapping  --------------------------------------
        okUH(0)             <= i_clk;
        okUH(1)             <= internal_if.hi_drive;
        okUH(4 downto 2)    <= internal_if.hi_cmd;
        internal_if.hi_datain <= okUHU;
        internal_if.hi_busy   <= okHU(0);
        okUHU               <= internal_if.hi_dataout when (internal_if.hi_drive = '1') else (others => 'Z');
        --end loop;
    end okHost_driver;

    -----------------------------------------------------------------------
    -- FrontPanelReset
    -----------------------------------------------------------------------
    procedure FrontPanelReset(signal i_clk : in std_logic; variable front_panel_conf : inout t_front_panel_conf; signal internal_if : inout t_internal_if) is
        variable i        : integer := 0;
        variable msg_line : line;
    begin
        for i in 31 downto 0 loop
            front_panel_conf.WireIns(i)   := (others => '0');
            front_panel_conf.WireOuts(i)  := (others => '0');
            front_panel_conf.Triggered(i) := (others => '0');
        end loop;
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd <= DReset;
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd <= DNOP;
        wait until (internal_if.hi_busy = '0');
    end procedure FrontPanelReset;

    -----------------------------------------------------------------------
    -- init_front_panel_record
    -----------------------------------------------------------------------
    impure function init_front_panel_conf(
         BlockDelayStates : in integer := 5; -- REQUIRED: # of clocks between blocks of pipe data
         ReadyCheckDelay  : in integer := 5; -- REQUIRED: # of clocks before block transfer before host interface checks for ready (0-255)
         PostReadyDelay   : in integer := 5; -- REQUIRED: # of clocks after ready is asserted and check that the block transfer begins (0-255)
         pipeInSize       : in integer := 1024; -- REQUIRED: byte (must be even) length of default PipeIn; Integer 0-2^32
         pipeOutSize      : in integer := 1024; -- REQUIRED: byte (must be even) length of default PipeOut; Integer 0-2^32
         registerSetSize  : in integer := 32 -- Size of array for register set commands.
    ) return t_front_panel_conf is

        variable result : t_front_panel_conf(
            pipeIn(0 to pipeInSize - 1),
            pipeOut(0 to pipeOutSize - 1),
            WireIns(0 to 31),
            WireOuts(0 to 31),
            Triggered(0 to 31),
            u32Address(0 to registerSetSize - 1),
            u32Data(0 to registerSetSize - 1)
        );

    begin
        result.PostReadyDelay   := PostReadyDelay;
        result.ReadyCheckDelay  := ReadyCheckDelay;
        result.BlockDelayStates := BlockDelayStates;
        result.pipeIn := (others => (others => '0'));
        result.pipeOut := (others => (others => '0'));
        result.WireIns := (others => (others => '0'));
        result.WireOuts := (others => (others => '0'));
        result.Triggered := (others => (others => '0'));

        return result;
    end function;

    -----------------------------------------------------------------------
    -- init_internal_if
    -----------------------------------------------------------------------
    impure function init_internal_if(
         dummy : in integer
    ) return t_internal_if is

        variable result : t_internal_if;
    begin
        result.hi_drive   := '0';
        result.hi_cmd  := (others => '0');
        result.hi_busy := '0';
        result.hi_datain := (others => '0');
        result.hi_dataout := (others => '0');

        return result;
    end function;

    -----------------------------------------------------------------------
    -- SetWireInValue
    -----------------------------------------------------------------------
    procedure SetWireInValue(
        ep                   : in std_logic_vector(7 downto 0);
        val                  : in std_logic_vector(31 downto 0);
        mask                 : in std_logic_vector(31 downto 0);
        variable front_panel_conf : inout t_front_panel_conf
    ) is

        variable tmp_slv32 : std_logic_vector(31 downto 0);
        variable tmpI      : integer;
    begin
        tmpI                      := to_integer(unsigned(ep));
        tmp_slv32                 := front_panel_conf.WireIns(tmpI) and (not mask);
        front_panel_conf.WireIns(tmpI) := (tmp_slv32 or (val and mask));
    end procedure SetWireInValue;

    -----------------------------------------------------------------------
    -- GetWireOutValue
    -----------------------------------------------------------------------
    impure function GetWireOutValue(
        ep          : std_logic_vector;
        front_panel_conf : in t_front_panel_conf)
    return std_logic_vector is

        variable tmp_slv32 : std_logic_vector(31 downto 0);
        variable tmpI      : integer;
    begin
        tmpI      := to_integer(unsigned(ep));
        tmp_slv32 := front_panel_conf.WireOuts(tmpI - 16#20#);
        return (tmp_slv32);
    end GetWireOutValue;

    -----------------------------------------------------------------------
    -- IsTriggered
    -----------------------------------------------------------------------
    impure function IsTriggered(
        ep          : std_logic_vector;
        mask        : std_logic_vector(31 downto 0);
        front_panel_conf : t_front_panel_conf
    ) return boolean is

        variable tmp_slv32 : std_logic_vector(front_panel_conf.Triggered(0)'range);
        variable tmpI      : integer;
        variable msg_line  : line;
    begin
        tmpI      := to_integer(unsigned(ep));
        tmp_slv32 := (front_panel_conf.Triggered(tmpI - 16#60#) and mask);

        if (tmp_slv32 >= std_logic_vector(to_unsigned(0, tmp_slv32'length))) then
            if (tmp_slv32 = std_logic_vector(to_unsigned(0, tmp_slv32'length))) then
                return FALSE;
            else
                return TRUE;
            end if;
        else
            write(msg_line, STRING'("***FRONTPANEL ERROR: IsTriggered mask 0x"));
            hwrite(msg_line, mask);
            write(msg_line, STRING'(" covers unused Triggers"));
            writeline(output, msg_line);
            return FALSE;
        end if;
    end IsTriggered;

    -----------------------------------------------------------------------
    -- UpdateWireIns
    -----------------------------------------------------------------------
    procedure UpdateWireIns(signal   i_clk   : in std_logic;
                            variable front_panel_conf : inout t_front_panel_conf;
                            signal   internal_if   : inout t_internal_if) is
        variable i : integer := 0;
    begin
        wait until (rising_edge(i_clk));
        wait for 12 ps;
        internal_if.hi_cmd   <= DWires;
        wait until (rising_edge(i_clk));
        wait for 12 ps;
        internal_if.hi_cmd   <= DUpdateWireIns;
        wait until (rising_edge(i_clk));
        wait for 12 ps;
        internal_if.hi_drive <= '1';
        wait until (rising_edge(i_clk));
        wait for 12 ps;
        internal_if.hi_cmd   <= DNOP;
        for i in 0 to 31 loop
            internal_if.hi_dataout <= front_panel_conf.WireIns(i);
            wait until (rising_edge(i_clk));
        wait for 12 ps;
        end loop;
        wait until (internal_if.hi_busy = '0');
    end procedure UpdateWireIns;

    -----------------------------------------------------------------------
    -- UpdateWireOuts
    -----------------------------------------------------------------------
    procedure UpdateWireOuts(
        signal   i_clk   : in std_logic;
        variable front_panel_conf : inout t_front_panel_conf;
        signal   internal_if   : inout t_internal_if
    ) is
        variable i : integer := 0;
    begin
        wait until (rising_edge(i_clk));
        wait for 12 ps;
        internal_if.hi_cmd   <= DWires;
        wait until (rising_edge(i_clk));
        wait for 12 ps;
        internal_if.hi_cmd   <= DUpdateWireOuts;
        wait until (rising_edge(i_clk));
        wait for 12 ps;
        wait until (rising_edge(i_clk));
        wait for 12 ps;
        internal_if.hi_cmd   <= DNOP;
        wait until (rising_edge(i_clk));
        wait for 12 ps;
        internal_if.hi_drive <= '0';
        wait until (rising_edge(i_clk));
        wait for 12 ps;
        wait until (rising_edge(i_clk));
        wait for 12 ps;
        for i in 0 to 31 loop
            wait until (rising_edge(i_clk));
            wait for 12 ps;
            front_panel_conf.WireOuts(i) := internal_if.hi_datain;
        end loop;
        wait until (internal_if.hi_busy = '0');
    end procedure UpdateWireOuts;

    -----------------------------------------------------------------------
    -- ActivateTriggerIn
    -----------------------------------------------------------------------
    procedure ActivateTriggerIn(
        signal i_clk : in std_logic;
        ep               : in std_logic_vector(7 downto 0);
        bit              : in integer;
        signal internal_if : inout t_internal_if) is

        variable tmp_slv5 : std_logic_vector(4 downto 0);
        variable c_ONE    : unsigned(31 downto 0) := x"00000001";
    begin
        tmp_slv5             := std_logic_vector(to_unsigned(bit, tmp_slv5'length));
        wait until (rising_edge(i_clk));
        wait for 12 ps;
        internal_if.hi_cmd     <= DTriggers;
        wait until (rising_edge(i_clk));
        wait for 12 ps;
        internal_if.hi_cmd     <= DActivateTriggerIn;
        wait until (rising_edge(i_clk));
        wait for 12 ps;
        internal_if.hi_drive   <= '1';
        internal_if.hi_dataout <= (x"000000" & ep);
        wait until (rising_edge(i_clk));
        wait for 12 ps;
        --hi_dataout <= SHL(x"00000001", tmp_slv5); 
        internal_if.hi_dataout <= std_logic_vector(c_ONE sll to_integer(unsigned(tmp_slv5))); -- TODO
        internal_if.hi_cmd     <= DNOP;
        wait until (rising_edge(i_clk));
        wait for 12 ps;
        internal_if.hi_dataout <= x"00000000";
        wait until (internal_if.hi_busy = '0');
    end procedure ActivateTriggerIn;

    -----------------------------------------------------------------------
    -- UpdateTriggerOuts
    -----------------------------------------------------------------------
    procedure UpdateTriggerOuts(
        signal   i_clk   : in std_logic;
        variable front_panel_conf : inout t_front_panel_conf;
        signal   internal_if   : inout t_internal_if
    ) is
    begin
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd   <= DTriggers;
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd   <= DUpdateTriggerOuts;
        wait until (rising_edge(i_clk));
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd   <= DNOP;
        wait until (rising_edge(i_clk));
        internal_if.hi_drive <= '0';
        wait until (rising_edge(i_clk));
        wait until (rising_edge(i_clk));
        wait until (rising_edge(i_clk));

        for i in 0 to (UPDATE_TO_READOUT_CLOCKS - 1) loop
            wait until (rising_edge(i_clk));
        end loop;

        for i in 0 to 31 loop
            wait until (rising_edge(i_clk));
            front_panel_conf.Triggered(i) := internal_if.hi_datain;
        end loop;
        wait until (internal_if.hi_busy = '0');
    end procedure UpdateTriggerOuts;

    -----------------------------------------------------------------------
    -- WriteToPipeIn
    -----------------------------------------------------------------------
    procedure WriteToPipeIn(
        signal   i_clk   : in std_logic;
        ep                   : in std_logic_vector(7 downto 0);
        length               : in integer;
        variable front_panel_conf : inout t_front_panel_conf;
        signal   internal_if   : inout t_internal_if) is

        variable len, i, j, k, blockSize : integer;
        variable tmp_slv8                : std_logic_vector(7 downto 0);
        variable tmp_slv32               : std_logic_vector(31 downto 0);
    begin
        len                  := (length / 4);
        j                    := 0;
        k                    := 0;
        blockSize            := 1024;
        tmp_slv8             := std_logic_vector(to_unsigned(front_panel_conf.BlockDelayStates, tmp_slv8'length));
        tmp_slv32            := std_logic_vector(to_unsigned(len, tmp_slv32'length));
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd     <= DPipes;
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd     <= DWriteToPipeIn;
        wait until (rising_edge(i_clk));
        internal_if.hi_drive   <= '1';
        internal_if.hi_dataout <= (x"0000" & tmp_slv8 & ep);
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd     <= DNOP;
        internal_if.hi_dataout <= tmp_slv32;
        for i in 0 to len - 1 loop
            wait until (rising_edge(i_clk));
            internal_if.hi_dataout(7 downto 0)   <= front_panel_conf.pipeIn(i * 4);
            internal_if.hi_dataout(15 downto 8)  <= front_panel_conf.pipeIn((i * 4) + 1);
            internal_if.hi_dataout(23 downto 16) <= front_panel_conf.pipeIn((i * 4) + 2);
            internal_if.hi_dataout(31 downto 24) <= front_panel_conf.pipeIn((i * 4) + 3);
            j                                  := j + 4;
            if (j = blockSize) then
                for k in 0 to front_panel_conf.BlockDelayStates - 1 loop
                    wait until (rising_edge(i_clk));
                end loop;
                j := 0;
            end if;
        end loop;
        wait until (internal_if.hi_busy = '0');
    end procedure WriteToPipeIn;

    -----------------------------------------------------------------------
    -- ReadFromPipeOut
    -----------------------------------------------------------------------
    procedure ReadFromPipeOut(
        signal   i_clk   : in std_logic;
        ep                   : in std_logic_vector(7 downto 0);
        length               : in integer;
        variable front_panel_conf : inout t_front_panel_conf;
        signal   internal_if   : inout t_internal_if
    ) is

        variable len, i, j, k, blockSize : integer;
        variable tmp_slv8                : std_logic_vector(7 downto 0);
        variable tmp_slv32               : std_logic_vector(31 downto 0);
    begin
        len                  := (length / 4);
        j                    := 0;
        blockSize            := 1024;
        tmp_slv8             := std_logic_vector(to_unsigned(front_panel_conf.BlockDelayStates, tmp_slv8'length));
        tmp_slv32            := std_logic_vector(to_unsigned(len, tmp_slv32'length));
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd     <= DPipes;
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd     <= DReadFromPipeOut;
        wait until (rising_edge(i_clk));
        internal_if.hi_drive   <= '1';
        internal_if.hi_dataout <= (x"0000" & tmp_slv8 & ep);
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd     <= DNOP;
        internal_if.hi_dataout <= tmp_slv32;
        wait until (rising_edge(i_clk));
        internal_if.hi_drive   <= '0';
        for i in 0 to len - 1 loop
            wait until (rising_edge(i_clk));
            front_panel_conf.pipeOut(i * 4)       := internal_if.hi_datain(7 downto 0);
            front_panel_conf.pipeOut((i * 4) + 1) := internal_if.hi_datain(15 downto 8);
            front_panel_conf.pipeOut((i * 4) + 2) := internal_if.hi_datain(23 downto 16);
            front_panel_conf.pipeOut((i * 4) + 3) := internal_if.hi_datain(31 downto 24);
            j                                := j + 4;
            if (j = blockSize) then
                for k in 0 to front_panel_conf.BlockDelayStates - 1 loop
                    wait until (rising_edge(i_clk));
                end loop;
                j := 0;
            end if;
        end loop;
        wait until (internal_if.hi_busy = '0');
    end procedure ReadFromPipeOut;

    -----------------------------------------------------------------------
    -- WriteToBlockPipeIn
    -----------------------------------------------------------------------
    procedure WriteToBlockPipeIn(
        signal   i_clk   : in std_logic;
        ep                   : in std_logic_vector(7 downto 0);
        blockLength          : in integer;
        length               : in integer;
        variable front_panel_conf : inout t_front_panel_conf;
        signal   internal_if   : inout t_internal_if) is

        variable len, i, j, k, blockSize, blockNum : integer;
        variable tmp_slv8                          : std_logic_vector(7 downto 0);
        variable tmp_slv16                         : std_logic_vector(15 downto 0);
        variable tmp_slv32                         : std_logic_vector(31 downto 0);
    begin
        len       := (length / 4);
        blockSize := (blockLength / 4);
        j         := 0;
        k         := 0;
        blockNum  := (len / blockSize);
        tmp_slv8  := std_logic_vector(to_unsigned(front_panel_conf.BlockDelayStates, tmp_slv8'length));
        tmp_slv16 := std_logic_vector(to_unsigned(blockSize, tmp_slv16'length));
        tmp_slv32 := std_logic_vector(to_unsigned(len, tmp_slv32'length));

        wait until (rising_edge(i_clk));
        internal_if.hi_cmd       <= DPipes;
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd       <= DWriteToBlockPipeIn;
        wait until (rising_edge(i_clk));
        internal_if.hi_drive     <= '1';
        internal_if.hi_dataout   <= (x"0000" & tmp_slv8 & ep);
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd       <= DNOP;
        internal_if.hi_dataout   <= tmp_slv32;
        wait until (rising_edge(i_clk));
        internal_if.hi_dataout   <= x"0000" & tmp_slv16;
        wait until (rising_edge(i_clk));
        tmp_slv16(15 downto 8) := std_logic_vector(to_unsigned(front_panel_conf.PostReadyDelay, 8));
        tmp_slv16(7 downto 0)  := std_logic_vector(to_unsigned(front_panel_conf.ReadyCheckDelay, 8));
        internal_if.hi_dataout   <= x"0000" & tmp_slv16;
        for i in 1 to blockNum loop
            while (internal_if.hi_busy = '1') loop
                wait until (rising_edge(i_clk));
            end loop;
            while (internal_if.hi_busy = '0') loop
                wait until (rising_edge(i_clk));
            end loop;
            wait until (rising_edge(i_clk));
            wait until (rising_edge(i_clk));
            for j in 1 to blockSize loop
                internal_if.hi_dataout(7 downto 0)   <= front_panel_conf.pipeIn(k);
                internal_if.hi_dataout(15 downto 8)  <= front_panel_conf.pipeIn(k + 1);
                internal_if.hi_dataout(23 downto 16) <= front_panel_conf.pipeIn(k + 2);
                internal_if.hi_dataout(31 downto 24) <= front_panel_conf.pipeIn(k + 3);
                wait until (rising_edge(i_clk));
                k                                  := k + 4;
            end loop;
            for j in 1 to front_panel_conf.BlockDelayStates loop
                wait until (rising_edge(i_clk));
            end loop;
        end loop;
        wait until (internal_if.hi_busy = '0');
    end procedure WriteToBlockPipeIn;

    -----------------------------------------------------------------------
    -- ReadFromBlockPipeOut
    -----------------------------------------------------------------------
    procedure ReadFromBlockPipeOut(
        signal   i_clk   : in std_logic;
        ep                   : in std_logic_vector(7 downto 0);
        blockLength          : in integer;
        length               : in integer;
        variable front_panel_conf : inout t_front_panel_conf;
        signal   internal_if   : inout t_internal_if) is

        variable len, i, j, k, blockSize, blockNum : integer;
        variable tmp_slv8                          : std_logic_vector(7 downto 0);
        variable tmp_slv16                         : std_logic_vector(15 downto 0);
        variable tmp_slv32                         : std_logic_vector(31 downto 0);
    begin
        len                    := (length / 4);
        blockSize              := (blockLength / 4);
        j                      := 0;
        k                      := 0;
        blockNum               := (len / blockSize);
        tmp_slv8               := std_logic_vector(to_unsigned(front_panel_conf.BlockDelayStates, tmp_slv8'length));
        tmp_slv16              := std_logic_vector(to_unsigned(blockSize, tmp_slv16'length));
        tmp_slv32              := std_logic_vector(to_unsigned(len, tmp_slv32'length));
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd       <= DPipes;
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd       <= DReadFromBlockPipeOut;
        wait until (rising_edge(i_clk));
        internal_if.hi_drive     <= '1';
        internal_if.hi_dataout   <= (x"0000" & tmp_slv8 & ep);
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd       <= DNOP;
        internal_if.hi_dataout   <= tmp_slv32;
        wait until (rising_edge(i_clk));
        internal_if.hi_dataout   <= x"0000" & tmp_slv16;
        wait until (rising_edge(i_clk));
        tmp_slv16(15 downto 8) := std_logic_vector(to_unsigned(front_panel_conf.PostReadyDelay, 8));
        tmp_slv16(7 downto 0)  := std_logic_vector(to_unsigned(front_panel_conf.ReadyCheckDelay, 8));
        internal_if.hi_dataout   <= x"0000" & tmp_slv16;
        wait until (rising_edge(i_clk));
        internal_if.hi_drive     <= '0';
        for i in 1 to blockNum loop
            while (internal_if.hi_busy = '1') loop
                wait until (rising_edge(i_clk));
            end loop;
            while (internal_if.hi_busy = '0') loop
                wait until (rising_edge(i_clk));
            end loop;
            wait until (rising_edge(i_clk));
            wait until (rising_edge(i_clk));
            for j in 1 to blockSize loop
                front_panel_conf.pipeOut(k)     := internal_if.hi_datain(7 downto 0);
                front_panel_conf.pipeOut(k + 1) := internal_if.hi_datain(15 downto 8);
                front_panel_conf.pipeOut(k + 2) := internal_if.hi_datain(23 downto 16);
                front_panel_conf.pipeOut(k + 3) := internal_if.hi_datain(31 downto 24);
                wait until (rising_edge(i_clk));
                k                          := k + 4;
            end loop;
            for j in 1 to front_panel_conf.BlockDelayStates loop
                wait until (rising_edge(i_clk));
            end loop;
        end loop;
        wait until (internal_if.hi_busy = '0');
    end procedure ReadFromBlockPipeOut;

    -----------------------------------------------------------------------
    -- WriteRegister
    -----------------------------------------------------------------------
    procedure WriteRegister(
        signal i_clk : in std_logic;
        address          : in std_logic_vector(31 downto 0);
        data             : in std_logic_vector(31 downto 0);
        signal internal_if : inout t_internal_if) is
    begin
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd     <= DRegisters;
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd     <= DWriteRegister;
        wait until (rising_edge(i_clk));
        internal_if.hi_drive   <= '1';
        internal_if.hi_cmd     <= DNOP;
        wait until (rising_edge(i_clk));
        internal_if.hi_dataout <= address;
        wait until (rising_edge(i_clk));
        internal_if.hi_dataout <= data;
        wait until (internal_if.hi_busy = '0');
        internal_if.hi_drive   <= '0';
    end procedure WriteRegister;

    -----------------------------------------------------------------------
    -- ReadRegister
    -----------------------------------------------------------------------
    procedure ReadRegister(
        signal i_clk : in std_logic;
        address          : in std_logic_vector(31 downto 0);
        data             : out std_logic_vector(31 downto 0);
        signal internal_if : inout t_internal_if) is
    begin
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd     <= DRegisters;
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd     <= DReadRegister;
        wait until (rising_edge(i_clk));
        internal_if.hi_drive   <= '1';
        internal_if.hi_cmd     <= DNOP;
        wait until (rising_edge(i_clk));
        internal_if.hi_dataout <= address;
        wait until (rising_edge(i_clk));
        internal_if.hi_drive   <= '0';
        wait until (rising_edge(i_clk));
        wait until (rising_edge(i_clk));
        data                 := internal_if.hi_datain;
        wait until (internal_if.hi_busy = '0');
    end procedure ReadRegister;

    -----------------------------------------------------------------------
    -- WriteRegisterSet
    -----------------------------------------------------------------------
    procedure WriteRegisterSet(
        signal   i_clk   : in std_logic;
        variable front_panel_conf : inout t_front_panel_conf;
        signal   internal_if   : inout t_internal_if) is
        variable i            : integer;
        variable u32Count_int : integer;
    begin
        u32Count_int         := to_integer(unsigned(front_panel_conf.u32Count));
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd     <= DRegisters;
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd     <= DWriteRegisterSet;
        wait until (rising_edge(i_clk));
        internal_if.hi_drive   <= '1';
        internal_if.hi_cmd     <= DNOP;
        wait until (rising_edge(i_clk));
        internal_if.hi_dataout <= front_panel_conf.u32Count;
        for i in 1 to u32Count_int loop
            wait until (rising_edge(i_clk));
            internal_if.hi_dataout <= front_panel_conf.u32Address(i - 1);
            wait until (rising_edge(i_clk));
            internal_if.hi_dataout <= front_panel_conf.u32Data(i - 1);
            wait until (rising_edge(i_clk));
            wait until (rising_edge(i_clk));
        end loop;
        wait until (internal_if.hi_busy = '0');
        internal_if.hi_drive   <= '0';
    end procedure WriteRegisterSet;

    -----------------------------------------------------------------------
    -- ReadRegisterSet
    -----------------------------------------------------------------------
    procedure ReadRegisterSet(
        signal   i_clk   : in std_logic;
        variable front_panel_conf : inout t_front_panel_conf;
        signal   internal_if   : inout t_internal_if
    ) is
        variable i            : integer;
        variable u32Count_int : integer;
    begin
        u32Count_int         := to_integer(unsigned(front_panel_conf.u32Count));
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd     <= DRegisters;
        wait until (rising_edge(i_clk));
        internal_if.hi_cmd     <= DReadRegisterSet;
        wait until (rising_edge(i_clk));
        internal_if.hi_drive   <= '1';
        internal_if.hi_cmd     <= DNOP;
        wait until (rising_edge(i_clk));
        internal_if.hi_dataout <= front_panel_conf.u32Count;
        for i in 1 to u32Count_int loop
            wait until (rising_edge(i_clk));
            internal_if.hi_dataout       <= front_panel_conf.u32Address(i - 1);
            wait until (rising_edge(i_clk));
            internal_if.hi_drive         <= '0';
            wait until (rising_edge(i_clk));
            wait until (rising_edge(i_clk));
            front_panel_conf.u32Data(i - 1) := internal_if.hi_datain;
            internal_if.hi_drive         <= '1';
        end loop;
        wait until (internal_if.hi_busy = '0');
    end procedure ReadRegisterSet;

end;
