-- -------------------------------------------------------------------------------------------------------------
--                              Copyright (C) 2022-2030 Ken-ji de la Rosa, IRAP Toulouse.
-- -------------------------------------------------------------------------------------------------------------
--                              This file is part of the ATHENA X-IFU DRE Focal Plane Assembly simulator.
--
--                              fpasim-fw is free software: you can redistribute it and/or modify
--                              it under the terms of the GNU General Public License as published by
--                              the Free Software Foundation, either version 3 of the License, or
--                              (at your option) any later version.
--
--                              This program is distributed in the hope that it will be useful,
--                              but WITHOUT ANY WARRANTY; without even the implied warranty of
--                              MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--                              GNU General Public License for more details.
--
--                              You should have received a copy of the GNU General Public License
--                              along with this program.  If not, see <https://www.gnu.org/licenses/>.
-- -------------------------------------------------------------------------------------------------------------
--    email                   kenji.delarosa@alten.com
--!   @file                   dac_frame_generator.vhd 
-- -------------------------------------------------------------------------------------------------------------
--    Automatic Generation    No
--    Code Rules Reference    SOC of design and VHDL handbook for VLSI development, CNES Edition (v2.1)
-- -------------------------------------------------------------------------------------------------------------
--!   @details                
--
-- This module generates flags to tags
--  . the first frame sample after the startup
--
--  Example0: continuous data valid signal
--  i_data_valid |   1   1   1   1   1   1   1   1   1   1   1   1   0   |   
--  o_sof        |   x   1   0   0   0   0   0   0   0   0   0   0   0   |
--  o_data_valid |   x   1   1   1   1   1   1   1   1   1   1   1   1   |
--
--  Example1: non-continuous data valid signal
--  g_frame_size |                   4                                                           |
--  i_data_valid |   1   0   1   0   1   0   1   0   1   0   1   0   1   0   1   0   1    0   1  |   
--  o_sof        |   1   0   0   0   0   0   0   0   0   0   0   0   0   0   0   0   0    0   0  |
--  o_data_valid |   1   0   1   0   1   0   1   0   1   0   1   0   1   0   1   0   1    0   1  |
--
-- -------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.pkg_utils;

entity dac_frame_generator is
  generic (
     g_DATA_WIDTH : integer := 16
     );
  port(
    i_clk        : in std_logic;        -- clock signal
    i_rst        : in std_logic;        -- reset signal
    ---------------------------------------------------------------------
    -- input
    ---------------------------------------------------------------------
    i_data_valid : in std_logic;        -- input valid sample
    i_data       : in std_logic_vector(g_DATA_WIDTH - 1 downto 0); -- input data

    ---------------------------------------------------------------------
    -- output
    ---------------------------------------------------------------------
    o_sof        : out std_logic;       -- first sample of the frame
    o_data_valid : out std_logic;        -- output valid sample
    o_data       : out std_logic_vector(g_DATA_WIDTH - 1  downto 0)
    );
end entity dac_frame_generator;

architecture RTL of dac_frame_generator is

  type t_state is (E_RST, E_WAIT, E_RUN);
  signal sm_state_r1   : t_state := E_RST;
  signal sm_state_next : t_state;

  signal sof_next : std_logic;
  signal sof_r1   : std_logic := '0';

  signal data_valid_next : std_logic;
  signal data_valid_r1   : std_logic := '0';

  signal data_r1 : std_logic_vector(o_data'range) := (others => '0');


begin

  -------------------------------------------------------------------
  -- fsm
  -------------------------------------------------------------------
  p_decode_state : process(sm_state_r1, i_data_valid) is
  begin
    sof_next        <= '0';
    data_valid_next <= '0';
    case sm_state_r1 is
      when E_RST =>
        sm_state_next <= E_WAIT;
      when E_WAIT =>
        if i_data_valid = '1' then
          sof_next        <= '1';
          data_valid_next <= i_data_valid;
          sm_state_next   <= E_RUN;
        else
          sm_state_next <= E_WAIT;
        end if;
      when E_RUN =>  -- @suppress "Dead state 'E_RUN': state does not have outgoing transitions"
        if i_data_valid = '1' then
          data_valid_next <= i_data_valid;
          sm_state_next   <= E_RUN;
        else
          sm_state_next <= E_RUN;
        end if;

      when others =>  -- @suppress "Case statement contains all choices explicitly. You can safely remove the redundant 'others'"
        sm_state_next <= E_RST;
    end case;
  end process p_decode_state;

  p_state : process(i_clk) is
  begin
    if rising_edge(i_clk) then
      if i_rst = '1' then
        sm_state_r1 <= E_RST;
      else
        sm_state_r1 <= sm_state_next;
      end if;
      sof_r1        <= sof_next;
      data_valid_r1 <= data_valid_next;

     -- pipe
     data_r1 <= i_data;

    end if;
  end process p_state;

  -------------------------------------------------------------------
  -- output
  -------------------------------------------------------------------
  o_sof        <= sof_r1;
  o_data_valid <= data_valid_r1;
  o_data       <= data_r1;

end architecture RTL;
